module multi
#(parameter radix = 78)
(
	input [radix-1:0] a,
	input [radix-1:0] b,
    input clk,
	output [42:0] res_0,
	output [42:0] res_1,
	output [42:0] res_2,
	output [42:0] res_3,
	output [42:0] res_4,
	output [42:0] res_5,
    output [42:0] res_6,
	output [42:0] res_7,
	output [42:0] res_8,
	output [42:0] res_9,
	output [42:0] res_10,
	output [42:0] res_11,
    output [42:0] res_12,
	output [42:0] res_13,
	output [42:0] res_14
);
    
    // this part needs to be changed based on the radix
	wire [25:0] wire_a [2:0];
	wire [16:0] wire_b [4:0];
    wire [42:0] result [14:0];
	assign wire_a[0] = a[25:0];
	assign wire_a[1] = a[51:26];
    assign wire_a[2] = a[77:52];
	assign wire_b[0] = b[16:0];
	assign wire_b[1] = b[33:17];
	assign wire_b[2] = b[50:34];
    assign wire_b[3] = b[67:51];
	assign wire_b[4] = {7'b0,b[77:68]};

    /***************************************/
    assign res_0 = result[0];
    assign res_1 = result[1];
    assign res_2 = result[2];
    assign res_3 = result[3];
    assign res_4 = result[4];
    assign res_5 = result[5];
    assign res_6 = result[6];
    assign res_7 = result[7];
    assign res_8 = result[8];
    assign res_9 = result[9];
    assign res_10 = result[10];
    assign res_11 = result[11];
    assign res_12 = result[12];
    assign res_13 = result[13];
    assign res_14 = result[14];

     genvar i;
     generate
         for(i=0;i<5;i=i+1) begin: dsp_generate
             dsp_macro_0 inst_dsp_0(
                 .CLK(clk),
                 .A(wire_a[0]),
                 .B(wire_b[i]),
                 .P({result[i]}));

             dsp_macro_0 inst_dsp_1(
                 .CLK(clk),
                 .A(wire_a[1]),
                 .B(wire_b[i]),
                 .P({result[i+5]}));

             dsp_macro_0 inst_dsp_2(
                 .CLK(clk),
                 .A(wire_a[2]),
                 .B(wire_b[i]),
                 .P({result[i+10]}));
         end
     endgenerate
    
	//original code(DSP slice usage is not well-scheduled)
    // assign res_0 = wire_a[0]*wire_b[0];
    // assign res_1 = wire_a[0]*wire_b[1];
    // assign res_2 = wire_a[0]*wire_b[2];
    // assign res_3 = wire_a[0]*wire_b[3];
    // assign res_4 = wire_a[0]*wire_b[4];
    // assign res_5 = wire_a[1]*wire_b[0];
    // assign res_6 = wire_a[1]*wire_b[1];
    // assign res_7 = wire_a[1]*wire_b[2];
    // assign res_8 = wire_a[1]*wire_b[3];
    // assign res_9 = wire_a[1]*wire_b[4];
    // assign res_10 = wire_a[2]*wire_b[0];
    // assign res_11 = wire_a[2]*wire_b[1];
    // assign res_12 = wire_a[2]*wire_b[2];
    // assign res_13 = wire_a[2]*wire_b[3];
    // assign res_14 = wire_a[2]*wire_b[4];
endmodule